VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM32
  CLASS BLOCK ;
  FOREIGN RAM32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 401.580 BY 136.000 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 399.580 17.720 401.580 18.320 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 399.580 29.960 401.580 30.560 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 399.580 42.200 401.580 42.800 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 399.580 54.440 401.580 55.040 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 399.580 66.680 401.580 67.280 ;
    END
  END A0[4]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 399.580 78.920 401.580 79.520 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 134.000 8.190 136.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 134.000 132.390 136.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 134.000 144.810 136.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 134.000 157.230 136.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 134.000 169.650 136.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 134.000 182.070 136.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 134.000 194.490 136.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 134.000 206.910 136.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 134.000 219.330 136.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 134.000 231.750 136.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 134.000 244.170 136.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 134.000 20.610 136.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 134.000 256.590 136.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 134.000 269.010 136.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 134.000 281.430 136.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 134.000 293.850 136.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 134.000 306.270 136.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 134.000 318.690 136.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 134.000 331.110 136.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 134.000 343.530 136.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 134.000 355.950 136.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 134.000 368.370 136.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 134.000 33.030 136.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 134.000 380.790 136.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 134.000 393.210 136.000 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 134.000 45.450 136.000 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 134.000 57.870 136.000 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 134.000 70.290 136.000 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 134.000 82.710 136.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 134.000 95.130 136.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 134.000 107.550 136.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 134.000 119.970 136.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 2.000 4.720 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 2.000 45.520 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 2.000 49.600 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 2.000 53.680 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 2.000 57.760 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 2.000 61.840 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 2.000 65.920 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 2.000 70.000 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 2.000 74.080 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 2.000 78.160 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 2.000 82.240 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 2.000 8.800 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 2.000 86.320 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 2.000 90.400 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 2.000 94.480 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 2.000 98.560 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 2.000 102.640 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 2.000 106.720 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 2.000 110.800 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 2.000 114.880 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 2.000 118.960 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 2.000 123.040 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 2.000 12.880 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 2.000 127.120 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 2.000 131.200 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 2.000 16.960 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 2.000 21.040 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 2.000 25.120 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 2.000 29.200 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 2.000 33.280 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 2.000 37.360 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 2.000 41.440 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 399.580 5.480 401.580 6.080 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.080 2.480 96.680 133.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.680 2.480 250.280 133.520 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 133.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.880 2.480 173.480 133.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.480 2.480 327.080 133.520 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 399.580 91.160 401.580 91.760 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 399.580 103.400 401.580 104.000 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 399.580 115.640 401.580 116.240 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 399.580 127.880 401.580 128.480 ;
    END
  END WE0[3]
  OBS
      LAYER li1 ;
        RECT 2.760 2.635 398.820 133.365 ;
      LAYER met1 ;
        RECT 2.460 0.040 398.820 135.960 ;
      LAYER met2 ;
        RECT 3.310 133.720 7.630 135.990 ;
        RECT 8.470 133.720 20.050 135.990 ;
        RECT 20.890 133.720 32.470 135.990 ;
        RECT 33.310 133.720 44.890 135.990 ;
        RECT 45.730 133.720 57.310 135.990 ;
        RECT 58.150 133.720 69.730 135.990 ;
        RECT 70.570 133.720 82.150 135.990 ;
        RECT 82.990 133.720 94.570 135.990 ;
        RECT 95.410 133.720 106.990 135.990 ;
        RECT 107.830 133.720 119.410 135.990 ;
        RECT 120.250 133.720 131.830 135.990 ;
        RECT 132.670 133.720 144.250 135.990 ;
        RECT 145.090 133.720 156.670 135.990 ;
        RECT 157.510 133.720 169.090 135.990 ;
        RECT 169.930 133.720 181.510 135.990 ;
        RECT 182.350 133.720 193.930 135.990 ;
        RECT 194.770 133.720 206.350 135.990 ;
        RECT 207.190 133.720 218.770 135.990 ;
        RECT 219.610 133.720 231.190 135.990 ;
        RECT 232.030 133.720 243.610 135.990 ;
        RECT 244.450 133.720 256.030 135.990 ;
        RECT 256.870 133.720 268.450 135.990 ;
        RECT 269.290 133.720 280.870 135.990 ;
        RECT 281.710 133.720 293.290 135.990 ;
        RECT 294.130 133.720 305.710 135.990 ;
        RECT 306.550 133.720 318.130 135.990 ;
        RECT 318.970 133.720 330.550 135.990 ;
        RECT 331.390 133.720 342.970 135.990 ;
        RECT 343.810 133.720 355.390 135.990 ;
        RECT 356.230 133.720 367.810 135.990 ;
        RECT 368.650 133.720 380.230 135.990 ;
        RECT 381.070 133.720 392.650 135.990 ;
        RECT 393.490 133.720 398.270 135.990 ;
        RECT 3.310 0.010 398.270 133.720 ;
      LAYER met3 ;
        RECT 2.000 131.600 399.580 133.445 ;
        RECT 2.400 130.200 399.580 131.600 ;
        RECT 2.000 128.880 399.580 130.200 ;
        RECT 2.000 127.520 399.180 128.880 ;
        RECT 2.400 127.480 399.180 127.520 ;
        RECT 2.400 126.120 399.580 127.480 ;
        RECT 2.000 123.440 399.580 126.120 ;
        RECT 2.400 122.040 399.580 123.440 ;
        RECT 2.000 119.360 399.580 122.040 ;
        RECT 2.400 117.960 399.580 119.360 ;
        RECT 2.000 116.640 399.580 117.960 ;
        RECT 2.000 115.280 399.180 116.640 ;
        RECT 2.400 115.240 399.180 115.280 ;
        RECT 2.400 113.880 399.580 115.240 ;
        RECT 2.000 111.200 399.580 113.880 ;
        RECT 2.400 109.800 399.580 111.200 ;
        RECT 2.000 107.120 399.580 109.800 ;
        RECT 2.400 105.720 399.580 107.120 ;
        RECT 2.000 104.400 399.580 105.720 ;
        RECT 2.000 103.040 399.180 104.400 ;
        RECT 2.400 103.000 399.180 103.040 ;
        RECT 2.400 101.640 399.580 103.000 ;
        RECT 2.000 98.960 399.580 101.640 ;
        RECT 2.400 97.560 399.580 98.960 ;
        RECT 2.000 94.880 399.580 97.560 ;
        RECT 2.400 93.480 399.580 94.880 ;
        RECT 2.000 92.160 399.580 93.480 ;
        RECT 2.000 90.800 399.180 92.160 ;
        RECT 2.400 90.760 399.180 90.800 ;
        RECT 2.400 89.400 399.580 90.760 ;
        RECT 2.000 86.720 399.580 89.400 ;
        RECT 2.400 85.320 399.580 86.720 ;
        RECT 2.000 82.640 399.580 85.320 ;
        RECT 2.400 81.240 399.580 82.640 ;
        RECT 2.000 79.920 399.580 81.240 ;
        RECT 2.000 78.560 399.180 79.920 ;
        RECT 2.400 78.520 399.180 78.560 ;
        RECT 2.400 77.160 399.580 78.520 ;
        RECT 2.000 74.480 399.580 77.160 ;
        RECT 2.400 73.080 399.580 74.480 ;
        RECT 2.000 70.400 399.580 73.080 ;
        RECT 2.400 69.000 399.580 70.400 ;
        RECT 2.000 67.680 399.580 69.000 ;
        RECT 2.000 66.320 399.180 67.680 ;
        RECT 2.400 66.280 399.180 66.320 ;
        RECT 2.400 64.920 399.580 66.280 ;
        RECT 2.000 62.240 399.580 64.920 ;
        RECT 2.400 60.840 399.580 62.240 ;
        RECT 2.000 58.160 399.580 60.840 ;
        RECT 2.400 56.760 399.580 58.160 ;
        RECT 2.000 55.440 399.580 56.760 ;
        RECT 2.000 54.080 399.180 55.440 ;
        RECT 2.400 54.040 399.180 54.080 ;
        RECT 2.400 52.680 399.580 54.040 ;
        RECT 2.000 50.000 399.580 52.680 ;
        RECT 2.400 48.600 399.580 50.000 ;
        RECT 2.000 45.920 399.580 48.600 ;
        RECT 2.400 44.520 399.580 45.920 ;
        RECT 2.000 43.200 399.580 44.520 ;
        RECT 2.000 41.840 399.180 43.200 ;
        RECT 2.400 41.800 399.180 41.840 ;
        RECT 2.400 40.440 399.580 41.800 ;
        RECT 2.000 37.760 399.580 40.440 ;
        RECT 2.400 36.360 399.580 37.760 ;
        RECT 2.000 33.680 399.580 36.360 ;
        RECT 2.400 32.280 399.580 33.680 ;
        RECT 2.000 30.960 399.580 32.280 ;
        RECT 2.000 29.600 399.180 30.960 ;
        RECT 2.400 29.560 399.180 29.600 ;
        RECT 2.400 28.200 399.580 29.560 ;
        RECT 2.000 25.520 399.580 28.200 ;
        RECT 2.400 24.120 399.580 25.520 ;
        RECT 2.000 21.440 399.580 24.120 ;
        RECT 2.400 20.040 399.580 21.440 ;
        RECT 2.000 18.720 399.580 20.040 ;
        RECT 2.000 17.360 399.180 18.720 ;
        RECT 2.400 17.320 399.180 17.360 ;
        RECT 2.400 15.960 399.580 17.320 ;
        RECT 2.000 13.280 399.580 15.960 ;
        RECT 2.400 11.880 399.580 13.280 ;
        RECT 2.000 9.200 399.580 11.880 ;
        RECT 2.400 7.800 399.580 9.200 ;
        RECT 2.000 6.480 399.580 7.800 ;
        RECT 2.000 5.120 399.180 6.480 ;
        RECT 2.400 5.080 399.180 5.120 ;
        RECT 2.400 3.720 399.580 5.080 ;
        RECT 2.000 0.855 399.580 3.720 ;
      LAYER met4 ;
        RECT 391.295 19.895 391.625 78.705 ;
  END
END RAM32
END LIBRARY

